module IF(
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	input [31:0]PC_OUT,
	input FLUSH,
	input PC_WRITE,
	input BRANCH,
	output [31:0]PC_4,
	output [31:0]instruction);

//TODO

endmodule