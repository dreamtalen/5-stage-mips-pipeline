module MEM(
	input clk,
	input rst_n,
	input [31:0]EX_MEM_aluOut,
	input [31:0]EX_MEM_writeData,
	input memWrite,
	input memRead,
	output [31:0]memReadData);

//TODO

endmodule